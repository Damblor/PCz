CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
769 79 2305 832
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
769 79 2305 832
177209362 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 170 406 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 189 360 0 1 11
0 10
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
12 SPDT Switch~
164 196 455 0 3 11
0 4 3 4
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3618 0 0
0
0
7 Pulser~
4 123 503 0 10 12
0 11 12 4 13 0 0 5 5 5
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6153 0 0
0
0
14 Logic Display~
6 251 198 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 227 200 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 212 200 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 190 198 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
9 2-In AND~
219 344 296 0 3 22
0 6 7 5
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3549 0 0
0
0
6 74LS90
107 219 302 0 10 21
0 10 10 5 5 4 8 9 6 7
8
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U1
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
14
3 3 4 0 0 8320 2 3 4 0 0 4
179 459
161 459
161 494
147 494
1 2 3 0 0 8320 0 1 3 0 0 6
182 406
187 406
187 446
174 446
174 451
179 451
1 5 4 0 0 8320 0 3 10 0 0 3
213 455
237 455
237 334
3 4 5 0 0 8320 0 9 10 0 0 4
342 319
342 342
219 342
219 328
1 0 6 0 0 8320 0 9 0 0 10 3
351 274
351 241
210 241
2 0 7 0 0 8320 0 9 0 0 9 3
333 274
333 251
227 251
6 0 8 0 0 12416 0 10 0 0 8 5
246 334
246 338
261 338
261 248
246 248
10 1 8 0 0 0 0 10 5 0 0 4
246 264
246 224
251 224
251 216
1 9 7 0 0 0 0 6 10 0 0 4
227 218
227 256
228 256
228 264
8 1 6 0 0 0 0 10 7 0 0 4
210 264
210 226
212 226
212 218
1 7 9 0 0 4224 0 8 10 0 0 4
190 216
190 256
192 256
192 264
1 1 10 0 0 4224 0 10 2 0 0 4
192 328
192 340
190 340
190 347
3 4 5 0 0 0 0 10 10 0 0 3
210 328
210 328
219 328
1 2 10 0 0 0 0 10 10 0 0 3
192 328
192 328
201 328
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
