CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
768 71 2304 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
768 71 2304 824
177209362 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 60 381 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 56 343 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 68 240 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
9 4-In AND~
219 571 188 0 5 22
0 6 5 4 3 10
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U6A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 542801386
65 0 0 0 2 1 6 0
1 U
6153 0 0
0
0
9 3-In AND~
219 437 182 0 4 22
0 6 5 4 7
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 5 0
1 U
5394 0 0
0
0
6 JK RN~
219 633 289 0 6 22
0 10 9 10 8 15 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U4A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 4 0
1 U
7734 0 0
0
0
12 Hex Display~
7 81 28 0 16 19
10 2 16 17 18 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
9914 0 0
0
0
12 Hex Display~
7 116 28 0 18 19
10 6 5 4 3 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3747 0 0
0
0
12 SPDT Switch~
164 83 339 0 10 11
0 9 9 14 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3549 0 0
0
0
7 Pulser~
4 33 293 0 10 12
0 19 20 21 9 0 0 5 5 2
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7931 0 0
0
0
9 2-In AND~
219 317 180 0 3 22
0 6 5 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9325 0 0
0
0
6 JK RN~
219 506 283 0 6 22
0 7 9 7 8 22 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
8903 0 0
0
0
6 JK RN~
219 370 281 0 6 22
0 11 9 11 8 23 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3834 0 0
0
0
6 JK RN~
219 254 284 0 6 22
0 6 9 6 8 24 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
3363 0 0
0
0
6 JK RN~
219 137 289 0 6 22
0 12 9 12 8 25 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
7668 0 0
0
0
42
1 5 2 0 0 4096 0 7 0 0 16 2
90 52
90 82
4 4 3 0 0 4096 0 8 0 0 16 2
107 52
107 82
3 3 4 0 0 4096 0 8 0 0 16 4
113 52
113 77
114 77
114 82
2 2 5 0 0 4096 0 8 0 0 16 2
119 52
119 82
1 1 6 0 0 4096 0 8 0 0 16 2
125 52
125 82
6 5 2 0 0 8320 0 6 0 0 16 3
657 272
667 272
667 82
0 4 3 0 0 8320 0 0 0 10 16 3
541 232
472 232
472 82
0 3 4 0 0 8320 0 0 0 23 16 3
405 231
349 231
349 82
0 2 5 0 0 8192 0 0 0 25 16 3
288 220
266 220
266 82
6 4 3 0 0 0 0 12 4 0 0 4
530 266
541 266
541 202
547 202
0 1 6 0 0 8320 0 0 4 12 0 5
405 160
405 162
539 162
539 175
547 175
0 1 6 0 0 0 0 0 5 32 0 5
289 171
289 160
405 160
405 173
413 173
1 0 7 0 0 4096 0 12 0 0 14 2
482 266
458 266
4 3 7 0 0 4224 0 5 12 0 0 3
458 182
458 284
482 284
1 0 6 0 0 0 0 0 0 16 32 2
211 82
211 171
5 0 1 0 0 4256 0 0 0 0 0 2
30 82
690 82
0 4 8 0 0 4096 0 0 6 31 0 3
506 381
633 381
633 320
0 2 9 0 0 4096 0 0 6 38 0 4
463 339
594 339
594 281
602 281
1 0 10 0 0 4096 0 6 0 0 20 2
609 272
596 272
5 3 10 0 0 8320 0 4 6 0 0 4
592 188
596 188
596 290
609 290
0 3 4 0 0 0 0 0 4 23 0 4
405 217
539 217
539 193
547 193
0 2 5 0 0 4224 0 0 4 25 0 4
288 208
532 208
532 184
547 184
6 3 4 0 0 0 0 13 5 0 0 4
394 264
405 264
405 191
413 191
0 2 5 0 0 0 0 0 5 25 0 4
288 201
405 201
405 182
413 182
6 2 5 0 0 0 0 14 11 0 0 4
278 267
288 267
288 189
293 189
1 0 11 0 0 4096 0 13 0 0 27 3
346 264
334 264
334 262
3 3 11 0 0 8320 0 11 13 0 0 6
338 180
342 180
342 245
334 245
334 282
346 282
4 0 8 0 0 0 0 15 0 0 31 4
137 320
137 376
138 376
138 381
4 0 8 0 0 0 0 14 0 0 31 2
254 315
254 381
4 0 8 0 0 0 0 13 0 0 31 2
370 312
370 381
1 4 8 0 0 4224 0 1 12 0 0 3
72 381
506 381
506 314
0 1 6 0 0 0 0 0 11 34 0 3
202 272
202 171
293 171
0 3 6 0 0 0 0 0 14 34 0 3
215 272
215 285
230 285
6 1 6 0 0 0 0 15 14 0 0 4
161 272
217 272
217 267
230 267
2 0 9 0 0 0 0 15 0 0 38 2
106 281
106 339
2 0 9 0 0 0 0 14 0 0 38 2
223 276
223 339
2 0 9 0 0 0 0 13 0 0 38 2
339 273
339 339
1 2 9 0 0 4224 0 9 12 0 0 4
100 339
464 339
464 275
475 275
1 0 12 0 0 4096 0 15 0 0 40 2
113 272
97 272
1 3 12 0 0 8320 0 3 15 0 0 4
80 240
97 240
97 290
113 290
4 2 9 0 0 4224 13 10 9 0 0 3
63 293
63 335
66 335
3 1 14 0 0 4224 0 9 2 0 0 2
66 343
68 343
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
