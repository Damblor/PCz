CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
42991634 0
0
6 Title:
5 Name:
0
0
0
37
13 Logic Switch~
5 248 339 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 121 469 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 871 67 0 1 11
0 17
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 679 62 0 1 11
0 16
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 515 61 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 356 69 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -23 8 -15
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 272 210 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9914 0 0
0
0
14 Logic Display~
6 944 487 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 847 495 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 746 494 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 636 495 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
12 D Flip-Flop~
219 888 549 0 4 9
0 4 7 31 3
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U9
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8903 0 0
0
0
12 D Flip-Flop~
219 789 549 0 4 9
0 5 7 32 4
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U8
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3834 0 0
0
0
12 D Flip-Flop~
219 685 549 0 4 9
0 6 7 33 5
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3363 0 0
0
0
12 D Flip-Flop~
219 576 549 0 4 9
0 2 7 34 6
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
7 Pulser~
4 115 405 0 10 12
0 35 36 7 37 0 0 5 5 4
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4718 0 0
0
0
12 SPDT Switch~
164 191 437 0 10 11
0 7 7 9 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3874 0 0
0
0
14 Logic Display~
6 908 329 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 719 333 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 552 330 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 399 333 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3750 0 0
0
0
9 Inverter~
13 899 97 0 2 22
0 17 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
8778 0 0
0
0
9 Inverter~
13 705 91 0 2 22
0 16 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
538 0 0
0
0
9 Inverter~
13 538 96 0 2 22
0 15 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
6843 0 0
0
0
9 Inverter~
13 382 101 0 2 22
0 14 21
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3136 0 0
0
0
9 2-In AND~
219 927 263 0 3 22
0 18 22 23
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
5950 0 0
0
0
9 2-In AND~
219 864 264 0 3 22
0 17 22 27
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5670 0 0
0
0
9 2-In AND~
219 736 262 0 3 22
0 19 22 24
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6828 0 0
0
0
9 2-In AND~
219 672 262 0 3 22
0 16 22 28
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6735 0 0
0
0
9 2-In AND~
219 568 262 0 3 22
0 20 22 25
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
8365 0 0
0
0
9 2-In AND~
219 508 263 0 3 22
0 15 22 29
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4132 0 0
0
0
9 2-In AND~
219 419 263 0 3 22
0 21 22 26
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4551 0 0
0
0
9 2-In AND~
219 349 265 0 3 22
0 14 22 30
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3635 0 0
0
0
5 4013~
219 862 386 0 6 22
0 27 11 7 23 38 2
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 2 2 0
1 U
3973 0 0
0
0
5 4013~
219 670 386 0 6 22
0 28 12 7 24 39 11
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 1 2 0
1 U
3851 0 0
0
0
5 4013~
219 506 386 0 6 22
0 29 13 7 25 40 12
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 2 1 0
1 U
8383 0 0
0
0
5 4013~
219 347 386 0 6 22
0 30 8 7 26 41 13
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 1 1 0
1 U
9334 0 0
0
0
54
0 1 2 0 0 8320 0 0 15 20 0 5
904 350
904 454
544 454
544 513
552 513
4 1 3 0 0 4224 0 12 8 0 0 3
912 513
944 513
944 505
1 0 4 0 0 0 0 9 0 0 10 2
847 513
847 513
1 0 5 0 0 4096 0 10 0 0 11 2
746 512
746 513
1 0 6 0 0 0 0 11 0 0 12 2
636 513
636 513
2 0 7 0 0 8192 0 15 0 0 9 3
552 531
548 531
548 546
2 0 7 0 0 0 0 14 0 0 9 3
661 531
657 531
657 546
2 0 7 0 0 0 0 13 0 0 9 3
765 531
761 531
761 546
0 2 7 0 0 8192 0 0 12 16 0 5
302 437
302 546
856 546
856 531
864 531
4 1 4 0 0 4224 0 13 12 0 0 2
813 513
864 513
4 1 5 0 0 4224 0 14 13 0 0 2
709 513
765 513
4 1 6 0 0 4224 0 15 14 0 0 2
600 513
661 513
3 0 7 0 0 0 0 37 0 0 16 3
323 368
313 368
313 437
3 0 7 0 0 0 0 36 0 0 16 3
482 368
473 368
473 437
3 0 7 0 0 0 0 35 0 0 16 3
646 368
643 368
643 437
1 3 7 0 0 4224 0 17 34 0 0 4
208 437
830 437
830 368
838 368
1 2 8 0 0 4224 0 1 37 0 0 4
260 339
315 339
315 350
323 350
3 1 9 0 0 4224 0 17 2 0 0 4
174 441
142 441
142 469
133 469
3 2 7 0 0 8320 10 16 17 0 0 4
139 396
166 396
166 433
174 433
1 6 2 0 0 128 0 18 34 0 0 3
908 347
908 350
886 350
1 0 11 0 0 4096 0 19 0 0 52 2
719 351
719 350
1 0 12 0 0 16 0 20 0 0 53 2
552 348
552 350
1 0 13 0 0 4096 0 21 0 0 54 2
399 351
399 350
1 0 14 0 0 4096 0 25 0 0 35 2
367 101
356 101
1 0 15 0 0 4096 0 24 0 0 34 2
523 96
515 96
1 0 16 0 0 4096 0 23 0 0 33 2
690 91
679 91
1 0 17 0 0 4096 0 22 0 0 32 2
884 97
871 97
1 2 18 0 0 4224 0 26 22 0 0 3
934 241
934 97
920 97
2 1 19 0 0 8320 0 23 28 0 0 3
726 91
743 91
743 240
1 2 20 0 0 4224 0 30 24 0 0 3
575 240
575 96
559 96
2 1 21 0 0 8320 0 25 32 0 0 3
403 101
426 101
426 241
1 1 17 0 0 4224 0 3 27 0 0 2
871 79
871 242
1 1 16 0 0 4224 0 29 4 0 0 2
679 240
679 74
1 1 15 0 0 4224 0 5 31 0 0 2
515 73
515 241
1 1 14 0 0 4224 0 6 33 0 0 2
356 81
356 243
2 0 22 0 0 4096 0 32 0 0 43 2
408 241
408 210
2 0 22 0 0 4096 0 33 0 0 43 2
338 243
338 210
2 0 22 0 0 0 0 31 0 0 43 2
497 241
497 210
2 0 22 0 0 0 0 30 0 0 43 2
557 240
557 210
2 0 22 0 0 0 0 29 0 0 43 4
661 240
661 215
662 215
662 210
2 0 22 0 0 0 0 28 0 0 43 2
725 240
725 210
2 0 22 0 0 0 0 27 0 0 43 2
853 242
853 210
1 2 22 0 0 4224 0 7 26 0 0 3
284 210
916 210
916 241
4 3 23 0 0 12416 0 34 26 0 0 4
862 392
862 396
925 396
925 286
4 3 24 0 0 12416 0 35 28 0 0 4
670 392
670 396
734 396
734 285
4 3 25 0 0 12416 0 36 30 0 0 4
506 392
506 396
566 396
566 285
4 3 26 0 0 12416 0 37 32 0 0 4
347 392
347 396
417 396
417 286
1 3 27 0 0 4224 0 34 27 0 0 2
862 329
862 287
3 1 28 0 0 4224 0 29 35 0 0 2
670 285
670 329
1 3 29 0 0 4224 0 36 31 0 0 2
506 329
506 286
3 1 30 0 0 4224 0 33 37 0 0 2
347 288
347 329
6 2 11 0 0 4224 0 35 34 0 0 4
694 350
849 350
849 350
838 350
6 2 12 0 0 4224 0 36 35 0 0 4
530 350
659 350
659 350
646 350
6 2 13 0 0 4224 0 37 36 0 0 2
371 350
482 350
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
