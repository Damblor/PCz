CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
769 79 1543 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
769 79 1543 831
177209362 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 413 357 0 1 11
0 8
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 381 355 0 1 11
0 9
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 151 363 0 1 11
0 14
0
0 0 21360 90
2 0V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 185 363 0 1 11
0 13
0
0 0 21360 90
2 0V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 70 436 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
7 Pulser~
4 67 504 0 10 12
0 17 18 19 4 0 0 5 5 2
7
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7734 0 0
0
0
12 SPDT Switch~
164 138 436 0 10 11
0 2 2 4 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
9914 0 0
0
0
14 Logic Display~
6 444 239 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 426 242 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 407 240 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 389 241 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
6 74LS90
107 416 293 0 10 21
0 9 9 8 8 6 7 12 11 10
7
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U1
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
6 74LS90
107 188 302 0 10 21
0 14 14 13 13 2 5 6 16 15
5
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U2
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3834 0 0
0
0
14 Logic Display~
6 161 247 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 179 250 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 197 248 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 214 249 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
22
1 5 2 0 0 8320 0 7 13 0 0 3
155 436
206 436
206 334
2 1 2 0 0 4224 3 7 5 0 0 4
121 432
91 432
91 436
82 436
4 3 4 0 0 8320 0 6 7 0 0 4
97 504
113 504
113 440
121 440
6 10 5 0 0 4224 0 13 13 0 0 2
215 334
215 264
7 5 6 0 0 8320 0 13 12 0 0 3
161 264
161 325
434 325
1 6 7 0 0 4224 0 8 12 0 0 3
444 257
444 325
443 325
4 0 8 0 0 4112 0 12 0 0 9 4
416 319
416 332
414 332
414 337
1 2 9 0 0 8336 0 2 12 0 0 4
382 342
382 333
398 333
398 319
3 1 8 0 0 4240 0 12 1 0 0 4
407 319
407 337
414 337
414 344
1 1 9 0 0 16 0 2 12 0 0 4
382 342
382 333
389 333
389 319
1 10 7 0 0 16 0 8 12 0 0 3
444 257
444 255
443 255
1 9 10 0 0 4240 0 9 12 0 0 3
426 260
426 255
425 255
1 8 11 0 0 4240 0 10 12 0 0 2
407 258
407 255
1 7 12 0 0 4240 0 11 12 0 0 2
389 259
389 255
1 4 13 0 0 12288 0 4 13 0 0 4
186 350
186 342
188 342
188 328
3 1 13 0 0 4224 0 13 4 0 0 4
179 328
179 343
186 343
186 350
2 1 14 0 0 8320 0 13 3 0 0 4
170 328
170 343
152 343
152 350
1 1 14 0 0 0 0 13 3 0 0 4
161 328
161 343
152 343
152 350
1 10 5 0 0 0 0 17 13 0 0 3
214 267
214 264
215 264
1 9 15 0 0 4224 0 16 13 0 0 2
197 266
197 264
1 8 16 0 0 4224 0 15 13 0 0 2
179 268
179 264
1 7 6 0 0 0 0 14 13 0 0 2
161 265
161 264
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
