CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
42991634 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 191 180 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 97 271 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 811 152 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 670 162 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 526 162 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 363 161 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
12 D Flip-Flop~
219 724 216 0 4 9
0 4 3 10 2
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U4
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
12 D Flip-Flop~
219 571 216 0 4 9
0 5 3 11 4
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3747 0 0
0
0
12 D Flip-Flop~
219 423 216 0 4 9
0 6 3 12 5
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
12 D Flip-Flop~
219 265 216 0 4 9
0 7 3 13 6
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
12 SPDT Switch~
164 167 239 0 10 11
0 3 3 8 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
9325 0 0
0
0
7 Pulser~
4 91 207 0 10 12
0 14 15 3 16 0 0 5 5 5
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8903 0 0
0
0
14
4 1 2 0 0 4224 0 7 3 0 0 3
748 180
811 180
811 170
2 0 3 0 0 8192 0 10 0 0 5 3
241 198
233 198
233 239
2 0 3 0 0 0 0 8 0 0 5 3
547 198
541 198
541 239
2 0 3 0 0 0 0 9 0 0 5 3
399 198
395 198
395 239
1 2 3 0 0 4224 0 11 7 0 0 4
184 239
692 239
692 198
700 198
1 0 4 0 0 0 0 4 0 0 9 2
670 180
670 180
1 0 5 0 0 0 0 5 0 0 10 2
526 180
526 180
1 0 6 0 0 4096 0 6 0 0 11 2
363 179
363 180
4 1 4 0 0 4224 0 8 7 0 0 2
595 180
700 180
4 1 5 0 0 4224 0 9 8 0 0 2
447 180
547 180
4 1 6 0 0 4224 0 10 9 0 0 2
289 180
399 180
1 1 7 0 0 4224 0 1 10 0 0 2
203 180
241 180
3 1 8 0 0 4224 0 11 2 0 0 4
150 243
118 243
118 271
109 271
3 2 3 0 0 8320 9 12 11 0 0 4
115 198
142 198
142 235
150 235
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
