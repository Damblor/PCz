CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
768 71 2304 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
768 71 2304 824
177209362 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 171 144 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 217 232 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 50 271 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 688 167 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 555 167 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 423 166 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 287 166 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
5 SCOPE
12 720 172 0 1 11
0 2
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 598 173 0 1 11
0 3
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 473 172 0 1 11
0 4
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 339 172 0 1 11
0 5
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9325 0 0
0
0
5 SCOPE
12 91 193 0 1 11
0 13
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8903 0 0
0
0
9 Inverter~
13 172 191 0 2 22
0 6 7
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3834 0 0
0
0
6 JK RN~
219 655 201 0 6 22
0 3 13 9 12 15 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
3363 0 0
0
0
6 JK RN~
219 514 201 0 6 22
0 4 13 10 12 9 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
7668 0 0
0
0
6 JK RN~
219 381 201 0 6 22
0 5 13 11 12 10 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
4718 0 0
0
0
6 JK RN~
219 248 201 0 6 22
0 6 13 7 12 11 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
3874 0 0
0
0
12 SPDT Switch~
164 120 248 0 10 11
0 13 13 14 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
6671 0 0
0
0
7 Pulser~
4 50 213 0 10 12
0 16 17 13 18 0 0 5 5 1
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3789 0 0
0
0
28
1 0 2 0 0 4096 0 4 0 0 8 2
688 185
688 184
1 0 3 0 0 4096 0 5 0 0 16 2
555 185
555 184
1 0 4 0 0 0 0 6 0 0 17 2
423 184
423 184
1 0 5 0 0 0 0 7 0 0 18 2
287 184
287 184
1 0 6 0 0 8192 0 1 0 0 7 3
183 144
188 144
188 169
2 3 7 0 0 8320 0 13 17 0 0 5
175 209
175 213
201 213
201 202
224 202
1 1 6 0 0 8336 0 13 17 0 0 5
175 173
175 169
205 169
205 184
224 184
6 1 2 0 0 4224 0 14 8 0 0 2
679 184
720 184
1 0 3 0 0 0 0 9 0 0 16 2
598 185
598 184
1 0 4 0 0 0 0 10 0 0 17 2
473 184
473 184
1 0 5 0 0 0 0 11 0 0 18 2
339 184
339 184
1 0 13 0 0 4096 8 12 0 0 28 2
91 205
91 204
5 3 9 0 0 4224 0 15 14 0 0 2
544 202
631 202
5 3 10 0 0 4224 0 16 15 0 0 2
411 202
490 202
5 3 11 0 0 4224 0 17 16 0 0 2
278 202
357 202
6 1 3 0 0 4224 0 15 14 0 0 2
538 184
631 184
6 1 4 0 0 4224 0 16 15 0 0 2
405 184
490 184
6 1 5 0 0 4224 0 17 16 0 0 2
272 184
357 184
4 4 12 0 0 4224 0 15 14 0 0 2
514 232
655 232
4 4 12 0 0 0 0 16 15 0 0 2
381 232
514 232
4 4 12 0 0 0 0 17 16 0 0 2
248 232
381 232
1 4 12 0 0 0 0 2 17 0 0 2
229 232
248 232
0 2 13 0 0 4224 0 0 14 24 0 4
471 248
613 248
613 193
624 193
0 2 13 0 0 0 0 0 15 25 0 4
342 248
471 248
471 193
483 193
0 2 13 0 0 0 0 0 16 26 0 4
209 248
342 248
342 193
350 193
1 2 13 0 0 0 0 18 17 0 0 4
137 248
209 248
209 193
217 193
3 1 14 0 0 4224 0 18 3 0 0 4
103 252
71 252
71 271
62 271
3 2 13 0 0 8320 8 19 18 0 0 4
74 204
95 204
95 244
103 244
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
