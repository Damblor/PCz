CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
769 79 1535 823
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
769 79 1535 823
177209362 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 22 375 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 116 259 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 99 260 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 82 259 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 64 258 0 1 11
0 6
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 48 259 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 31 257 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 13 256 0 1 11
0 3
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 360 206 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V12
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 337 206 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V11
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 314 207 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V10
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 290 207 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8903 0 0
0
0
14 Logic Display~
6 313 331 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
7 74LS151
20 203 327 0 14 29
0 9 8 7 6 5 4 3 2 13
12 11 10 14 15
0
0 0 13040 0
7 74LS151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3363 0 0
0
0
13
1 8 2 0 0 4224 0 1 14 0 0 4
34 375
163 375
163 363
171 363
1 7 3 0 0 8320 0 8 14 0 0 3
13 268
13 354
171 354
1 6 4 0 0 8320 0 7 14 0 0 3
31 269
31 345
171 345
5 1 5 0 0 4224 0 14 6 0 0 3
171 336
48 336
48 271
1 4 6 0 0 8320 0 5 14 0 0 3
64 270
64 327
171 327
3 1 7 0 0 4224 0 14 4 0 0 3
171 318
82 318
82 271
1 2 8 0 0 8320 0 3 14 0 0 3
99 272
99 309
171 309
1 1 9 0 0 4224 0 14 2 0 0 3
171 300
116 300
116 271
1 12 10 0 0 8320 0 9 14 0 0 5
360 218
360 315
249 315
249 327
235 327
11 1 11 0 0 8320 0 14 10 0 0 5
235 318
301 318
301 226
337 226
337 218
1 10 12 0 0 4224 0 11 14 0 0 3
314 219
314 309
235 309
9 1 13 0 0 8320 0 14 12 0 0 3
241 300
290 300
290 219
13 1 14 0 0 4224 0 14 13 0 0 3
235 354
313 354
313 349
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
