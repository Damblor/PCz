CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
177209362 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 217 199 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 97 271 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
5 SCOPE
12 774 291 0 1 11
0 2
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 684 125 0 1 11
0 3
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 517 125 0 1 11
0 4
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 341 126 0 1 11
0 5
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 207 228 0 1 11
0 6
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
14 Logic Display~
6 801 119 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 651 117 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 484 119 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 315 118 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
9 Inverter~
13 184 125 0 2 22
0 7 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
8903 0 0
0
0
9 Inverter~
13 449 303 0 2 22
0 2 9
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4D
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
3834 0 0
0
0
9 Inverter~
13 415 294 0 2 22
0 3 10
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
3363 0 0
0
0
9 Inverter~
13 381 285 0 2 22
0 4 11
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
7668 0 0
0
0
9 Inverter~
13 337 276 0 2 22
0 5 12
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
4718 0 0
0
0
10 4-In NAND~
219 269 290 0 5 22
0 9 10 11 12 7
0
0 0 624 180
6 74LS20
-21 -28 21 -20
3 U3A
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 3 0
1 U
3874 0 0
0
0
6 JK RN~
219 269 153 0 6 22
0 8 6 7 18 17 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
6671 0 0
0
0
6 JK RN~
219 439 153 0 6 22
0 5 6 17 18 16 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
3789 0 0
0
0
6 JK RN~
219 611 153 0 6 22
0 4 6 16 18 15 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
4871 0 0
0
0
6 JK RN~
219 768 153 0 6 22
0 3 6 15 18 19 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
3750 0 0
0
0
12 SPDT Switch~
164 167 239 0 3 11
0 6 14 6
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
8778 0 0
0
0
7 Pulser~
4 91 207 0 10 12
0 20 21 14 22 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
538 0 0
0
0
36
1 0 2 0 0 0 0 3 0 0 17 2
774 303
774 303
1 0 3 0 0 4096 0 4 0 0 28 2
684 137
684 136
1 0 4 0 0 4096 0 5 0 0 30 2
517 137
517 136
1 0 5 0 0 4096 0 6 0 0 32 2
341 138
341 136
1 0 6 0 0 4096 0 7 0 0 13 2
207 240
207 239
1 0 2 0 0 4096 0 8 0 0 17 2
801 137
801 136
1 0 3 0 0 0 0 9 0 0 28 2
651 135
651 136
1 0 4 0 0 0 0 10 0 0 30 2
484 137
484 136
1 0 5 0 0 0 0 11 0 0 32 2
315 136
315 136
0 2 6 0 0 4112 0 0 21 11 0 4
572 237
729 237
729 145
737 145
0 2 6 0 0 4224 0 0 20 12 0 4
390 237
572 237
572 145
580 145
2 0 6 0 0 0 0 19 0 0 13 5
408 145
390 145
390 238
233 238
233 239
1 2 6 0 0 0 0 22 18 0 0 4
184 239
235 239
235 145
238 145
5 0 7 0 0 8320 0 17 0 0 15 3
242 290
189 290
189 154
1 3 7 0 0 0 0 12 18 0 0 4
169 125
165 125
165 154
245 154
2 1 8 0 0 4224 0 12 18 0 0 4
205 125
230 125
230 136
245 136
1 6 2 0 0 4224 0 13 21 0 0 4
470 303
810 303
810 136
792 136
1 0 3 0 0 4224 0 14 0 0 28 3
436 294
716 294
716 136
1 0 4 0 0 4224 0 15 0 0 30 3
402 285
560 285
560 136
1 0 5 0 0 4224 0 16 0 0 32 2
358 276
358 136
2 1 9 0 0 4224 0 13 17 0 0 2
434 303
293 303
2 2 10 0 0 4224 0 14 17 0 0 2
400 294
293 294
2 3 11 0 0 4224 0 15 17 0 0 2
366 285
293 285
2 4 12 0 0 4224 0 16 17 0 0 2
322 276
293 276
3 1 6 0 0 4224 13 22 2 0 0 4
150 243
118 243
118 271
109 271
3 2 14 0 0 8320 0 23 22 0 0 4
115 198
142 198
142 235
150 235
5 3 15 0 0 4224 0 20 21 0 0 2
641 154
744 154
6 1 3 0 0 0 0 20 21 0 0 2
635 136
744 136
5 3 16 0 0 4224 0 19 20 0 0 2
469 154
587 154
6 1 4 0 0 0 0 19 20 0 0 2
463 136
587 136
5 3 17 0 0 4224 0 18 19 0 0 2
299 154
415 154
6 1 5 0 0 0 0 18 19 0 0 2
293 136
415 136
4 0 18 0 0 8192 0 21 0 0 34 3
768 184
768 197
611 197
4 0 18 0 0 8320 0 20 0 0 35 4
611 184
611 197
438 197
438 198
0 4 18 0 0 0 0 0 19 36 0 4
268 199
268 198
439 198
439 184
1 4 18 0 0 0 0 1 18 0 0 3
229 199
269 199
269 184
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
