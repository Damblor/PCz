CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
769 79 1535 823
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
769 79 1535 823
177209362 0
0
6 Title:
5 Name:
0
0
0
28
9 Inverter~
13 186 439 0 2 22
0 7 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
8953 0 0
0
0
9 Inverter~
13 187 527 0 2 22
0 8 3
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
4441 0 0
0
0
9 Inverter~
13 272 439 0 2 22
0 6 5
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3618 0 0
0
0
9 Inverter~
13 275 537 0 2 22
0 3 4
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
6153 0 0
0
0
10 3-In NAND~
219 402 406 0 4 22
0 3 6 2 9
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 4 0
1 U
5394 0 0
0
0
10 3-In NAND~
219 403 460 0 4 22
0 4 6 2 10
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 4 0
1 U
7734 0 0
0
0
10 3-In NAND~
219 405 511 0 4 22
0 5 3 2 11
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 3 0
1 U
9914 0 0
0
0
10 3-In NAND~
219 404 567 0 4 22
0 5 4 2 12
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 3 0
1 U
3747 0 0
0
0
14 Logic Display~
6 460 378 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 460 433 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 463 486 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 466 547 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
13 Logic Switch~
5 367 665 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21344 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 346 347 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3363 0 0
0
0
13 Logic Switch~
5 63 205 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7668 0 0
0
0
13 Logic Switch~
5 66 122 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4718 0 0
0
0
14 Logic Display~
6 445 229 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 442 168 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 439 115 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 439 60 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
10 3-In NAND~
219 383 249 0 4 22
0 5 4 2 12
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
3750 0 0
0
0
10 3-In NAND~
219 384 193 0 4 22
0 5 3 2 11
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 2 0
1 U
8778 0 0
0
0
10 3-In NAND~
219 382 142 0 4 22
0 4 6 2 10
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 2 0
1 U
538 0 0
0
0
10 3-In NAND~
219 381 88 0 4 22
0 3 6 2 9
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
6843 0 0
0
0
9 Inverter~
13 254 219 0 2 22
0 3 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3136 0 0
0
0
9 Inverter~
13 251 121 0 2 22
0 6 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
5950 0 0
0
0
9 Inverter~
13 166 209 0 2 22
0 8 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
5670 0 0
0
0
9 Inverter~
13 165 121 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6828 0 0
0
0
40
1 0 0 0 0 0 0 2 0 0 34 3
172 527
98 527
98 205
1 0 0 0 0 0 0 1 0 0 33 3
171 439
126 439
126 122
3 0 2 0 0 16 0 8 0 0 6 2
380 576
368 576
3 0 2 0 0 16 0 7 0 0 6 2
381 520
368 520
3 0 2 0 0 16 0 6 0 0 6 4
379 469
373 469
373 470
368 470
1 3 2 0 0 16 0 13 5 0 0 3
368 652
368 415
378 415
0 0 3 0 0 16 0 0 0 8 15 3
345 465
230 465
230 527
2 1 3 0 0 16 0 7 5 0 0 4
381 511
345 511
345 397
378 397
0 2 4 0 0 16 0 0 4 10 0 2
356 537
296 537
1 2 4 0 0 16 0 6 8 0 0 4
379 451
356 451
356 567
380 567
0 2 5 0 0 16 0 0 3 12 0 4
373 524
301 524
301 439
293 439
1 1 5 0 0 16 0 8 7 0 0 4
380 558
373 558
373 502
381 502
0 0 6 0 0 16 0 0 0 14 16 3
371 424
230 424
230 439
2 2 6 0 0 16 0 5 6 0 0 4
378 406
371 406
371 460
379 460
2 1 3 0 0 16 0 2 4 0 0 4
208 527
252 527
252 537
260 537
2 1 6 0 0 16 0 1 3 0 0 2
207 439
257 439
4 1 9 0 0 16 0 5 9 0 0 3
429 406
460 406
460 396
4 1 10 0 0 16 0 6 10 0 0 3
430 460
460 460
460 451
4 1 11 0 0 16 0 7 11 0 0 3
432 511
463 511
463 504
4 1 12 0 0 16 0 8 12 0 0 5
431 567
454 567
454 573
466 573
466 565
3 0 2 0 0 4096 0 21 0 0 24 2
359 258
347 258
3 0 2 0 0 4096 0 22 0 0 24 2
360 202
347 202
3 0 2 0 0 0 0 23 0 0 24 4
358 151
352 151
352 152
347 152
1 3 2 0 0 4224 0 14 24 0 0 3
347 334
347 97
357 97
0 0 3 0 0 4224 0 0 0 26 35 3
324 147
209 147
209 209
2 1 3 0 0 0 0 22 24 0 0 4
360 193
324 193
324 79
357 79
0 2 4 0 0 4096 0 0 25 28 0 2
335 219
275 219
1 2 4 0 0 8320 0 23 21 0 0 4
358 133
335 133
335 249
359 249
0 2 5 0 0 8320 0 0 26 30 0 4
352 206
280 206
280 121
272 121
1 1 5 0 0 0 0 21 22 0 0 4
359 240
352 240
352 184
360 184
0 0 6 0 0 4224 0 0 0 32 36 3
350 106
209 106
209 121
2 2 6 0 0 0 0 24 23 0 0 4
357 88
350 88
350 142
358 142
1 1 7 0 0 4224 0 16 28 0 0 4
78 122
142 122
142 121
150 121
1 1 8 0 0 4224 0 15 27 0 0 4
75 205
143 205
143 209
151 209
2 1 3 0 0 0 0 27 25 0 0 4
187 209
231 209
231 219
239 219
2 1 6 0 0 0 0 28 26 0 0 2
186 121
236 121
4 1 9 0 0 4224 0 24 20 0 0 3
408 88
439 88
439 78
4 1 10 0 0 4224 0 23 19 0 0 3
409 142
439 142
439 133
4 1 11 0 0 4224 0 22 18 0 0 3
411 193
442 193
442 186
4 1 12 0 0 4224 0 21 17 0 0 5
410 249
433 249
433 255
445 255
445 247
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
