CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
768 71 2304 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
768 71 2304 824
177209362 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 60 381 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 56 343 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 68 240 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 521 206 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 400 247 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 283 251 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 190 256 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
12 Hex Display~
7 116 28 0 18 19
10 5 4 3 2 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3747 0 0
0
0
12 SPDT Switch~
164 83 339 0 10 11
0 9 9 12 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3549 0 0
0
0
7 Pulser~
4 33 293 0 10 12
0 13 14 15 9 0 0 5 5 4
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7931 0 0
0
0
9 2-In AND~
219 434 188 0 3 22
0 8 3 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9325 0 0
0
0
9 2-In AND~
219 317 180 0 3 22
0 5 4 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8903 0 0
0
0
6 JK RN~
219 506 283 0 6 22
0 7 9 7 6 16 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
3834 0 0
0
0
6 JK RN~
219 370 281 0 6 22
0 8 9 8 6 17 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3363 0 0
0
0
6 JK RN~
219 254 284 0 6 22
0 5 9 5 6 18 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
7668 0 0
0
0
6 JK RN~
219 137 289 0 6 22
0 10 9 10 6 19 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
4718 0 0
0
0
35
4 4 2 0 0 4096 0 8 0 0 10 2
107 52
107 94
3 3 3 0 0 4096 0 8 0 0 10 2
113 52
113 94
2 2 4 0 0 4096 0 8 0 0 10 2
119 52
119 94
1 1 5 0 0 4096 0 8 0 0 10 2
125 52
125 94
1 0 2 0 0 0 0 4 0 0 6 2
521 224
521 222
4 6 2 0 0 4224 0 0 13 10 0 4
507 94
507 222
530 222
530 266
0 3 3 0 0 4224 0 0 0 20 10 2
404 199
404 94
0 2 4 0 0 4224 0 0 0 24 10 2
288 190
288 94
0 1 5 0 0 4224 0 0 0 27 10 2
172 272
172 94
4 0 1 0 0 4256 0 0 0 0 0 2
50 94
516 94
4 0 6 0 0 4096 0 16 0 0 14 4
137 320
137 376
138 376
138 381
4 0 6 0 0 4096 0 15 0 0 14 2
254 315
254 381
4 0 6 0 0 4096 0 14 0 0 14 2
370 312
370 381
1 4 6 0 0 4224 0 1 13 0 0 3
72 381
506 381
506 314
1 0 3 0 0 0 0 5 0 0 20 2
400 265
400 264
1 0 4 0 0 0 0 6 0 0 24 2
283 269
283 267
1 0 5 0 0 0 0 7 0 0 27 2
190 274
190 272
0 3 7 0 0 4096 0 0 13 19 0 3
467 266
467 284
482 284
3 1 7 0 0 8320 0 11 13 0 0 4
455 188
467 188
467 266
482 266
6 2 3 0 0 0 0 14 11 0 0 4
394 264
404 264
404 197
410 197
0 3 8 0 0 4096 0 0 14 22 0 3
331 264
331 282
346 282
0 1 8 0 0 4224 0 0 14 23 0 5
343 180
343 245
331 245
331 264
346 264
3 1 8 0 0 0 0 12 11 0 0 4
338 180
402 180
402 179
410 179
6 2 4 0 0 0 0 15 12 0 0 4
278 267
288 267
288 189
293 189
0 1 5 0 0 0 0 0 12 27 0 3
202 272
202 171
293 171
0 3 5 0 0 0 0 0 15 27 0 3
215 272
215 285
230 285
6 1 5 0 0 0 0 16 15 0 0 4
161 272
217 272
217 267
230 267
2 0 9 0 0 4096 0 16 0 0 31 2
106 281
106 339
2 0 9 0 0 4096 0 15 0 0 31 2
223 276
223 339
2 0 9 0 0 4096 0 14 0 0 31 2
339 273
339 339
1 2 9 0 0 4224 0 9 13 0 0 4
100 339
464 339
464 275
475 275
1 0 10 0 0 4096 0 16 0 0 33 2
113 272
97 272
1 3 10 0 0 8320 0 3 16 0 0 4
80 240
97 240
97 290
113 290
4 2 9 0 0 4224 11 10 9 0 0 3
63 293
63 335
66 335
3 1 12 0 0 4224 0 9 2 0 0 2
66 343
68 343
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
