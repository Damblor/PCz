CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
768 71 2304 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
768 71 2304 824
177209362 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 217 232 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 50 271 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
9 Inverter~
13 174 175 0 2 22
0 2 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
3618 0 0
0
0
9 Inverter~
13 415 318 0 2 22
0 4 8
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U3E
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
6153 0 0
0
0
9 Inverter~
13 379 309 0 2 22
0 5 9
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U3D
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
5394 0 0
0
0
9 Inverter~
13 346 300 0 2 22
0 6 10
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U3C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
7734 0 0
0
0
9 Inverter~
13 307 291 0 2 22
0 7 11
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U3B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
9914 0 0
0
0
10 4-In NAND~
219 239 305 0 5 22
0 8 9 10 11 2
0
0 0 624 180
6 74LS20
-21 -28 21 -20
3 U9A
-8 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 794459621
65 0 0 0 2 1 4 0
1 U
3747 0 0
0
0
14 Logic Display~
6 688 167 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 555 167 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 423 166 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 287 166 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
5 SCOPE
12 720 172 0 1 11
0 4
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3834 0 0
0
0
5 SCOPE
12 598 173 0 1 11
0 5
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3363 0 0
0
0
5 SCOPE
12 473 172 0 1 11
0 6
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7668 0 0
0
0
5 SCOPE
12 339 172 0 1 11
0 7
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4718 0 0
0
0
5 SCOPE
12 91 193 0 1 11
0 17
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3874 0 0
0
0
6 JK RN~
219 655 201 0 6 22
0 5 17 13 16 19 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
6671 0 0
0
0
6 JK RN~
219 514 201 0 6 22
0 6 17 14 16 13 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
3789 0 0
0
0
6 JK RN~
219 381 201 0 6 22
0 7 17 15 16 14 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
4871 0 0
0
0
6 JK RN~
219 248 201 0 6 22
0 3 17 2 16 15 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
3750 0 0
0
0
12 SPDT Switch~
164 120 248 0 10 11
0 17 17 18 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
8778 0 0
0
0
7 Pulser~
4 50 213 0 10 12
0 20 21 17 22 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
538 0 0
0
0
36
5 0 2 0 0 8320 0 8 0 0 2 3
212 305
169 305
169 202
1 3 2 0 0 0 0 3 21 0 0 4
159 175
155 175
155 202
224 202
2 1 3 0 0 12416 0 3 21 0 0 4
195 175
209 175
209 184
224 184
1 0 4 0 0 4224 0 4 0 0 16 3
436 318
701 318
701 184
1 0 5 0 0 4240 0 5 0 0 24 4
400 309
578 309
578 184
577 184
1 0 6 0 0 8320 0 6 0 0 25 3
367 300
440 300
440 184
1 0 7 0 0 8192 0 7 0 0 26 5
328 291
371 291
371 236
324 236
324 184
2 1 8 0 0 4224 0 4 8 0 0 2
400 318
263 318
2 2 9 0 0 4224 0 5 8 0 0 2
364 309
263 309
2 3 10 0 0 4224 0 6 8 0 0 2
331 300
263 300
2 4 11 0 0 4224 0 7 8 0 0 2
292 291
263 291
1 0 4 0 0 0 0 9 0 0 16 2
688 185
688 184
1 0 5 0 0 0 0 10 0 0 24 2
555 185
555 184
1 0 6 0 0 0 0 11 0 0 25 2
423 184
423 184
1 0 7 0 0 0 0 12 0 0 26 2
287 184
287 184
6 1 4 0 0 128 0 18 13 0 0 2
679 184
720 184
1 0 5 0 0 0 0 14 0 0 24 2
598 185
598 184
1 0 6 0 0 0 0 15 0 0 25 2
473 184
473 184
1 0 7 0 0 0 0 16 0 0 26 2
339 184
339 184
1 0 17 0 0 4096 12 17 0 0 36 2
91 205
91 204
5 3 13 0 0 4224 0 19 18 0 0 2
544 202
631 202
5 3 14 0 0 4224 0 20 19 0 0 2
411 202
490 202
5 3 15 0 0 4224 0 21 20 0 0 2
278 202
357 202
6 1 5 0 0 128 0 19 18 0 0 2
538 184
631 184
6 1 6 0 0 128 0 20 19 0 0 2
405 184
490 184
6 1 7 0 0 4224 0 21 20 0 0 2
272 184
357 184
4 4 16 0 0 4224 0 19 18 0 0 2
514 232
655 232
4 4 16 0 0 0 0 20 19 0 0 2
381 232
514 232
4 4 16 0 0 0 0 21 20 0 0 2
248 232
381 232
1 4 16 0 0 0 0 1 21 0 0 2
229 232
248 232
0 2 17 0 0 4224 0 0 18 32 0 4
471 248
613 248
613 193
624 193
0 2 17 0 0 0 0 0 19 33 0 4
342 248
471 248
471 193
483 193
0 2 17 0 0 0 0 0 20 34 0 4
209 248
342 248
342 193
350 193
1 2 17 0 0 0 0 22 21 0 0 4
137 248
209 248
209 193
217 193
3 1 18 0 0 4224 0 22 2 0 0 4
103 252
71 252
71 271
62 271
3 2 17 0 0 8320 12 23 22 0 0 4
74 204
95 204
95 244
103 244
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
