CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 636 1536 824
193986578 0
0
6 Title:
5 Name:
0
0
0
19
6 JK RN~
219 473 320 0 6 22
0 10 6 10 9 17 5
0
0 0 4704 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
8953 0 0
0
0
6 JK RN~
219 663 319 0 6 22
0 10 5 10 9 16 3
0
0 0 4704 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
4441 0 0
0
0
6 JK RN~
219 833 318 0 6 22
0 10 3 10 9 15 4
0
0 0 4704 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3618 0 0
0
0
6 JK RN~
219 1031 320 0 6 22
0 10 4 10 9 14 2
0
0 0 4704 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
6153 0 0
0
0
7 Pulser~
4 290 315 0 10 12
0 11 12 6 13 0 0 5 5 4
7
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
5394 0 0
0
0
12 Hex Display~
7 455 133 0 18 19
10 5 3 4 2 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
7734 0 0
0
0
5 SCOPE
12 364 296 0 1 11
0 6
0
0 0 57568 0
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 564 291 0 1 11
0 5
0
0 0 57568 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 744 290 0 1 11
0 3
0
0 0 57568 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 928 289 0 1 11
0 4
0
0 0 57568 0
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 1121 292 0 1 11
0 2
0
0 0 57568 0
3 TP5
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9325 0 0
0
0
12 SPDT Switch~
164 336 357 0 10 11
0 6 6 8 0 0 0 0 0 0
1
0
0 0 4704 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
8903 0 0
0
0
14 Logic Display~
6 528 285 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 894 284 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 713 285 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 1084 287 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
13 Logic Switch~
5 300 209 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3874 0 0
0
0
13 Logic Switch~
5 409 363 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6671 0 0
0
0
13 Logic Switch~
5 309 361 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3789 0 0
0
0
31
5 2 0 0 0 0 0 3 4 0 0 4
863 319
959 319
959 312
1000 312
5 2 0 0 0 0 0 2 3 0 0 4
693 320
772 320
772 310
802 310
5 2 0 0 0 0 0 1 2 0 0 4
503 321
599 321
599 311
632 311
1 0 2 0 0 16 0 16 0 0 12 2
1084 305
1084 304
1 0 3 0 0 16 0 15 0 0 14 2
713 303
713 302
1 0 4 0 0 16 0 14 0 0 13 2
894 302
894 301
1 0 5 0 0 16 0 13 0 0 15 2
528 303
528 303
0 1 5 0 0 16 0 0 6 15 0 4
506 303
506 188
464 188
464 157
0 2 3 0 0 16 0 0 6 14 0 4
694 302
694 184
458 184
458 157
0 3 4 0 0 16 0 0 6 13 0 4
871 301
871 178
452 178
452 157
0 4 2 0 0 16 0 0 6 12 0 4
1064 304
1064 172
446 172
446 157
6 1 2 0 0 16 0 4 11 0 0 3
1055 303
1055 304
1121 304
6 1 4 0 0 16 0 3 10 0 0 2
857 301
928 301
6 1 3 0 0 16 0 2 9 0 0 2
687 302
744 302
6 1 5 0 0 16 0 1 8 0 0 2
497 303
564 303
1 2 6 0 0 16 0 7 1 0 0 4
364 308
437 308
437 312
442 312
1 1 6 0 0 16 0 12 7 0 0 3
353 357
353 308
364 308
3 2 6 0 0 16 7 5 12 0 0 3
314 306
319 306
319 353
1 3 8 0 0 16 0 19 12 0 0 2
321 361
319 361
4 0 9 0 0 16 0 1 0 0 23 2
473 351
473 363
4 0 9 0 0 16 0 2 0 0 23 2
663 350
663 363
4 0 9 0 0 16 0 3 0 0 23 2
833 349
833 363
1 4 9 0 0 16 0 18 4 0 0 3
421 363
1031 363
1031 351
1 0 10 0 0 16 0 1 0 0 25 2
449 303
427 303
0 3 10 0 0 16 0 0 1 31 0 3
427 209
427 321
449 321
1 0 10 0 0 16 0 2 0 0 27 2
639 302
622 302
0 3 10 0 0 16 0 0 2 31 0 3
622 209
622 320
639 320
1 0 10 0 0 16 0 3 0 0 29 2
809 301
793 301
0 3 10 0 0 16 0 0 3 31 0 3
793 209
793 319
809 319
1 0 10 0 0 16 0 4 0 0 31 2
1007 303
983 303
1 3 10 0 0 16 0 17 4 0 0 4
312 209
983 209
983 321
1007 321
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
