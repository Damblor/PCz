CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
768 71 2304 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
768 71 2304 824
177209362 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 131 193 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 60 381 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 56 343 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 68 240 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6153 0 0
0
0
9 Inverter~
13 165 169 0 2 22
0 7 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
5394 0 0
0
0
9 3-In AND~
219 402 290 0 4 22
0 11 6 7 9
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 5 0
1 U
7734 0 0
0
0
9 3-In AND~
219 404 250 0 4 22
0 5 4 3 10
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 5 0
1 U
9914 0 0
0
0
8 2-In OR~
219 445 273 0 3 22
0 10 9 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3747 0 0
0
0
8 2-In OR~
219 257 278 0 3 22
0 15 16 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3549 0 0
0
0
9 2-In AND~
219 213 303 0 3 22
0 6 7 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7931 0 0
0
0
9 2-In AND~
219 213 259 0 3 22
0 5 4 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9325 0 0
0
0
12 Hex Display~
7 81 28 0 16 19
10 17 22 23 24 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
8903 0 0
0
0
12 Hex Display~
7 116 28 0 16 19
10 4 3 2 18 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3834 0 0
0
0
12 SPDT Switch~
164 83 339 0 10 11
0 8 8 21 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3363 0 0
0
0
7 Pulser~
4 33 293 0 10 12
0 25 26 27 8 0 0 5 5 1
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7668 0 0
0
0
6 JK RN~
219 511 276 0 6 22
0 13 8 13 12 28 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
4718 0 0
0
0
6 JK RN~
219 337 279 0 6 22
0 14 8 14 12 11 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
3874 0 0
0
0
6 JK RN~
219 137 289 0 6 22
0 19 8 19 12 6 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
6671 0 0
0
0
38
6 3 2 0 0 8320 0 16 0 0 34 3
535 259
545 259
545 82
0 2 3 0 0 12416 0 0 0 16 34 4
369 262
369 314
372 314
372 82
0 1 4 0 0 12288 0 0 0 26 34 4
173 272
173 183
191 183
191 82
0 2 4 0 0 8320 0 0 7 26 0 5
177 272
177 233
371 233
371 250
380 250
2 1 5 0 0 4224 0 5 7 0 0 4
186 169
356 169
356 241
380 241
1 2 5 0 0 0 0 11 5 0 0 6
189 250
185 250
185 183
191 183
191 169
186 169
0 2 6 0 0 12432 0 0 6 25 0 6
181 294
185 294
185 321
368 321
368 290
378 290
0 3 7 0 0 8320 0 0 6 9 0 5
167 312
167 333
372 333
372 299
378 299
1 2 7 0 0 0 0 1 10 0 0 4
143 193
167 193
167 312
189 312
1 1 7 0 0 0 0 1 5 0 0 6
143 193
148 193
148 183
145 183
145 169
150 169
0 2 8 0 0 8192 0 0 16 12 0 5
296 349
296 347
472 347
472 268
480 268
0 2 8 0 0 8320 0 0 17 13 0 5
103 339
103 349
298 349
298 271
306 271
1 2 8 0 0 0 0 14 18 0 0 6
100 339
104 339
104 324
101 324
101 281
106 281
2 4 9 0 0 8320 0 8 6 0 0 3
432 282
432 290
423 290
4 1 10 0 0 4224 0 7 8 0 0 3
425 250
425 264
432 264
3 6 3 0 0 0 0 7 17 0 0 4
380 259
375 259
375 262
361 262
5 1 11 0 0 12416 0 17 6 0 0 4
367 280
372 280
372 281
378 281
4 0 12 0 0 8192 0 16 0 0 27 3
511 307
511 376
337 376
1 3 13 0 0 4224 0 16 8 0 0 3
487 259
487 273
478 273
3 3 13 0 0 0 0 8 16 0 0 3
478 273
478 277
487 277
1 3 14 0 0 8320 0 17 9 0 0 4
313 262
298 262
298 278
290 278
3 3 14 0 0 0 0 9 17 0 0 4
290 278
298 278
298 280
313 280
3 1 15 0 0 4224 0 11 9 0 0 3
234 259
234 269
244 269
3 2 16 0 0 8320 0 10 9 0 0 4
234 303
238 303
238 287
244 287
5 1 6 0 0 0 0 18 10 0 0 4
167 290
181 290
181 294
189 294
6 2 4 0 0 0 0 18 11 0 0 4
161 272
181 272
181 268
189 268
4 0 12 0 0 8320 0 17 0 0 28 4
337 310
337 376
135 376
135 381
1 4 12 0 0 0 0 2 18 0 0 3
72 381
137 381
137 320
1 5 17 0 0 4224 0 12 0 0 34 2
90 52
90 82
4 4 18 0 0 4224 0 13 0 0 34 2
107 52
107 82
3 3 2 0 0 0 0 13 0 0 34 4
113 52
113 77
114 77
114 82
2 2 3 0 0 0 0 13 0 0 34 2
119 52
119 82
1 1 4 0 0 0 0 13 0 0 34 2
125 52
125 82
5 0 1 0 0 4256 0 0 0 0 0 2
30 82
690 82
1 0 19 0 0 4096 0 18 0 0 36 2
113 272
97 272
1 3 19 0 0 8320 0 4 18 0 0 4
80 240
97 240
97 290
113 290
4 2 8 0 0 4224 20 15 14 0 0 3
63 293
63 335
66 335
3 1 21 0 0 4224 0 14 3 0 0 2
66 343
68 343
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
