CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
42991634 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 248 339 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 121 469 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 871 67 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 679 62 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 515 61 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 356 69 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -23 8 -15
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 272 210 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
7 Pulser~
4 115 405 0 10 12
0 27 28 2 29 0 0 5 5 3
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3747 0 0
0
0
12 SPDT Switch~
164 191 437 0 10 11
0 2 2 4 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3549 0 0
0
0
14 Logic Display~
6 908 329 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 719 333 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 547 332 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 399 333 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
9 Inverter~
13 899 97 0 2 22
0 13 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
3363 0 0
0
0
9 Inverter~
13 705 91 0 2 22
0 12 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
7668 0 0
0
0
9 Inverter~
13 538 96 0 2 22
0 11 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
4718 0 0
0
0
9 Inverter~
13 382 101 0 2 22
0 10 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3874 0 0
0
0
9 2-In AND~
219 927 263 0 3 22
0 14 18 19
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
6671 0 0
0
0
9 2-In AND~
219 864 264 0 3 22
0 13 18 23
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3789 0 0
0
0
9 2-In AND~
219 736 262 0 3 22
0 15 18 20
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4871 0 0
0
0
9 2-In AND~
219 672 262 0 3 22
0 12 18 24
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3750 0 0
0
0
9 2-In AND~
219 568 262 0 3 22
0 16 18 21
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
8778 0 0
0
0
9 2-In AND~
219 508 263 0 3 22
0 11 18 25
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
538 0 0
0
0
9 2-In AND~
219 419 263 0 3 22
0 17 18 22
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6843 0 0
0
0
9 2-In AND~
219 349 265 0 3 22
0 10 18 26
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3136 0 0
0
0
5 4013~
219 862 386 0 6 22
0 23 7 2 19 30 6
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 2 2 0
1 U
5950 0 0
0
0
5 4013~
219 670 386 0 6 22
0 24 8 2 20 31 7
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 1 2 0
1 U
5670 0 0
0
0
5 4013~
219 506 386 0 6 22
0 25 9 2 21 32 8
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 2 1 0
1 U
6828 0 0
0
0
5 4013~
219 347 386 0 6 22
0 26 3 2 22 33 9
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
65 0 0 512 2 1 1 0
1 U
6735 0 0
0
0
42
3 0 2 0 0 8192 0 29 0 0 4 3
323 368
313 368
313 437
3 0 2 0 0 0 0 28 0 0 4 3
482 368
473 368
473 437
3 0 2 0 0 0 0 27 0 0 4 3
646 368
643 368
643 437
1 3 2 0 0 4224 0 9 26 0 0 4
208 437
830 437
830 368
838 368
1 2 3 0 0 4224 0 1 29 0 0 4
260 339
315 339
315 350
323 350
3 1 4 0 0 4240 0 9 2 0 0 4
174 441
142 441
142 469
133 469
3 2 2 0 0 8336 5 8 9 0 0 4
139 396
166 396
166 433
174 433
1 6 6 0 0 8320 0 10 26 0 0 3
908 347
908 350
886 350
1 0 7 0 0 4096 0 11 0 0 40 2
719 351
719 350
1 0 8 0 0 0 0 12 0 0 41 2
547 350
547 350
1 0 9 0 0 4096 0 13 0 0 42 2
399 351
399 350
1 0 10 0 0 4096 0 17 0 0 23 2
367 101
356 101
1 0 11 0 0 4096 0 16 0 0 22 2
523 96
515 96
1 0 12 0 0 4096 0 15 0 0 21 2
690 91
679 91
1 0 13 0 0 4096 0 14 0 0 20 2
884 97
871 97
1 2 14 0 0 4224 0 18 14 0 0 3
934 241
934 97
920 97
2 1 15 0 0 8320 0 15 20 0 0 3
726 91
743 91
743 240
1 2 16 0 0 4224 0 22 16 0 0 3
575 240
575 96
559 96
2 1 17 0 0 8320 0 17 24 0 0 3
403 101
426 101
426 241
1 1 13 0 0 4224 0 3 19 0 0 2
871 79
871 242
1 1 12 0 0 4224 0 21 4 0 0 2
679 240
679 74
1 1 11 0 0 4224 0 5 23 0 0 2
515 73
515 241
1 1 10 0 0 4224 0 6 25 0 0 2
356 81
356 243
2 0 18 0 0 4096 0 24 0 0 31 2
408 241
408 210
2 0 18 0 0 4096 0 25 0 0 31 2
338 243
338 210
2 0 18 0 0 0 0 23 0 0 31 2
497 241
497 210
2 0 18 0 0 0 0 22 0 0 31 2
557 240
557 210
2 0 18 0 0 0 0 21 0 0 31 4
661 240
661 215
662 215
662 210
2 0 18 0 0 0 0 20 0 0 31 2
725 240
725 210
2 0 18 0 0 0 0 19 0 0 31 2
853 242
853 210
1 2 18 0 0 4224 0 7 18 0 0 3
284 210
916 210
916 241
4 3 19 0 0 12416 0 26 18 0 0 4
862 392
862 396
925 396
925 286
4 3 20 0 0 12416 0 27 20 0 0 4
670 392
670 396
734 396
734 285
4 3 21 0 0 12416 0 28 22 0 0 4
506 392
506 396
566 396
566 285
4 3 22 0 0 12416 0 29 24 0 0 4
347 392
347 396
417 396
417 286
1 3 23 0 0 4224 0 26 19 0 0 2
862 329
862 287
3 1 24 0 0 4224 0 21 27 0 0 2
670 285
670 329
1 3 25 0 0 4224 0 28 23 0 0 2
506 329
506 286
3 1 26 0 0 4224 0 25 29 0 0 2
347 288
347 329
6 2 7 0 0 4224 0 27 26 0 0 4
694 350
849 350
849 350
838 350
6 2 8 0 0 4224 0 28 27 0 0 4
530 350
659 350
659 350
646 350
6 2 9 0 0 4224 0 29 28 0 0 2
371 350
482 350
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
