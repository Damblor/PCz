CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
177209362 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 300 209 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 309 361 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
9 Inverter~
13 1002 139 0 2 22
0 3 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3618 0 0
0
0
5 SCOPE
12 1118 128 0 1 11
0 2
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6153 0 0
0
0
9 3-In AND~
219 968 139 0 4 22
0 6 5 4 3
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
5394 0 0
0
0
6 JK RN~
219 473 320 0 6 22
0 11 8 11 2 12 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
7734 0 0
0
0
6 JK RN~
219 663 319 0 6 22
0 11 6 11 2 13 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
9914 0 0
0
0
6 JK RN~
219 833 318 0 6 22
0 11 5 11 2 14 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3747 0 0
0
0
6 JK RN~
219 1031 320 0 6 22
0 11 4 11 2 15 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
3549 0 0
0
0
7 Pulser~
4 290 315 0 10 12
0 16 17 8 18 0 0 5 5 5
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7931 0 0
0
0
12 Hex Display~
7 455 133 0 18 19
10 6 5 4 7 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9325 0 0
0
0
5 SCOPE
12 364 296 0 1 11
0 8
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
5 SCOPE
12 564 291 0 1 11
0 6
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
5 SCOPE
12 744 290 0 1 11
0 5
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
5 SCOPE
12 928 289 0 1 11
0 4
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7668 0 0
0
0
5 SCOPE
12 1121 292 0 1 11
0 7
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4718 0 0
0
0
12 SPDT Switch~
164 336 357 0 10 11
0 8 8 10 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3874 0 0
0
0
14 Logic Display~
6 528 285 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 894 284 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 713 285 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 1084 287 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
36
0 4 2 0 0 4096 0 0 6 12 0 3
663 371
473 371
473 351
2 1 2 0 0 0 0 3 4 0 0 3
1023 139
1023 140
1118 140
1 4 3 0 0 4224 0 3 5 0 0 2
987 139
989 139
0 3 4 0 0 4096 0 0 5 7 0 2
944 312
944 148
0 2 5 0 0 4096 0 0 5 8 0 3
773 310
773 139
944 139
0 1 6 0 0 8320 0 0 5 9 0 3
586 311
586 130
944 130
2 1 4 0 0 0 0 9 15 0 0 3
1000 312
928 312
928 301
2 1 5 0 0 0 0 8 14 0 0 3
802 310
744 310
744 302
2 1 6 0 0 0 0 7 13 0 0 3
632 311
564 311
564 303
4 1 2 0 0 12416 0 9 4 0 0 5
1031 351
1031 371
1144 371
1144 140
1118 140
4 0 2 0 0 0 0 8 0 0 10 3
833 349
833 371
1031 371
4 0 2 0 0 0 0 7 0 0 11 3
663 350
663 371
833 371
1 0 7 0 0 4096 0 21 0 0 21 2
1084 305
1084 304
1 0 5 0 0 0 0 20 0 0 23 2
713 303
713 302
1 0 4 0 0 0 0 19 0 0 22 2
894 302
894 301
1 0 6 0 0 0 0 18 0 0 24 2
528 303
528 303
0 1 6 0 0 128 0 0 11 24 0 4
506 303
506 188
464 188
464 157
0 2 5 0 0 8320 0 0 11 23 0 4
694 302
694 184
458 184
458 157
0 3 4 0 0 8320 0 0 11 22 0 4
871 301
871 178
452 178
452 157
0 4 7 0 0 8320 0 0 11 21 0 4
1064 304
1064 172
446 172
446 157
6 1 7 0 0 0 0 9 16 0 0 3
1055 303
1055 304
1121 304
6 1 4 0 0 0 0 8 15 0 0 2
857 301
928 301
6 1 5 0 0 0 0 7 14 0 0 2
687 302
744 302
6 1 6 0 0 0 0 6 13 0 0 2
497 303
564 303
1 2 8 0 0 4224 0 12 6 0 0 4
364 308
437 308
437 312
442 312
1 1 8 0 0 0 0 17 12 0 0 3
353 357
353 308
364 308
3 2 8 0 0 8320 9 10 17 0 0 3
314 306
319 306
319 353
1 3 10 0 0 4224 0 2 17 0 0 2
321 361
319 361
1 0 11 0 0 4096 0 6 0 0 30 2
449 303
427 303
0 3 11 0 0 4096 0 0 6 36 0 3
427 209
427 321
449 321
1 0 11 0 0 0 0 7 0 0 32 2
639 302
622 302
0 3 11 0 0 0 0 0 7 36 0 3
622 209
622 320
639 320
1 0 11 0 0 0 0 8 0 0 34 2
809 301
793 301
0 3 11 0 0 0 0 0 8 36 0 3
793 209
793 319
809 319
1 0 11 0 0 0 0 9 0 0 36 2
1007 303
983 303
1 3 11 0 0 4224 0 1 9 0 0 4
312 209
983 209
983 321
1007 321
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
