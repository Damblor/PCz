CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
177209362 0
0
6 Title:
5 Name:
0
0
0
32
13 Logic Switch~
5 402 538 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 300 209 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 409 363 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 309 361 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
9 Inverter~
13 861 469 0 2 22
0 17 18
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
5394 0 0
0
0
9 Inverter~
13 679 461 0 2 22
0 17 19
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11B
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
7734 0 0
0
0
9 Inverter~
13 489 473 0 2 22
0 17 20
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11A
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
9914 0 0
0
0
8 2-In OR~
219 960 469 0 3 22
0 12 11 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3747 0 0
0
0
8 2-In OR~
219 769 464 0 3 22
0 14 13 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3549 0 0
0
0
8 2-In OR~
219 597 474 0 3 22
0 16 15 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U10A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7931 0 0
0
0
9 2-In AND~
219 729 487 0 3 22
0 17 9 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9325 0 0
0
0
9 2-In AND~
219 729 434 0 3 22
0 6 19 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
8903 0 0
0
0
9 2-In AND~
219 906 499 0 3 22
0 17 8 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3834 0 0
0
0
9 2-In AND~
219 905 438 0 3 22
0 5 18 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3363 0 0
0
0
9 2-In AND~
219 545 501 0 3 22
0 17 10 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7668 0 0
0
0
9 2-In AND~
219 545 446 0 3 22
0 7 20 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4718 0 0
0
0
6 JK RN~
219 473 320 0 6 22
0 26 22 26 25 10 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
3874 0 0
0
0
6 JK RN~
219 663 319 0 6 22
0 26 4 26 25 9 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
6671 0 0
0
0
6 JK RN~
219 833 318 0 6 22
0 26 3 26 25 8 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
3789 0 0
0
0
6 JK RN~
219 1031 320 0 6 22
0 26 2 26 25 27 21
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
4871 0 0
0
0
7 Pulser~
4 290 315 0 10 12
0 28 29 23 30 0 0 5 5 2
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3750 0 0
0
0
12 Hex Display~
7 455 133 0 18 19
10 7 6 5 21 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8778 0 0
0
0
5 SCOPE
12 364 296 0 1 11
0 22
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
538 0 0
0
0
5 SCOPE
12 564 291 0 1 11
0 7
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6843 0 0
0
0
5 SCOPE
12 744 290 0 1 11
0 6
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3136 0 0
0
0
5 SCOPE
12 928 289 0 1 11
0 5
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5950 0 0
0
0
5 SCOPE
12 1121 292 0 1 11
0 21
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5670 0 0
0
0
12 SPDT Switch~
164 336 357 0 3 11
0 22 23 22
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6828 0 0
0
0
14 Logic Display~
6 528 285 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
14 Logic Display~
6 894 284 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8365 0 0
0
0
14 Logic Display~
6 713 285 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4132 0 0
0
0
14 Logic Display~
6 1084 287 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4551 0 0
0
0
52
3 2 2 0 0 4224 0 8 20 0 0 3
993 469
993 312
1000 312
3 2 3 0 0 4224 0 9 19 0 0 2
802 464
802 310
3 2 4 0 0 8320 0 10 18 0 0 3
630 474
632 474
632 311
0 1 5 0 0 8192 0 0 14 34 0 3
883 301
881 301
881 429
0 1 6 0 0 8192 0 0 12 35 0 3
706 302
705 302
705 425
0 1 7 0 0 4224 0 0 16 36 0 3
513 303
513 437
521 437
5 2 8 0 0 8320 0 19 13 0 0 4
863 319
876 319
876 508
882 508
5 2 9 0 0 8320 0 18 11 0 0 4
693 320
700 320
700 496
705 496
5 2 10 0 0 8320 0 17 15 0 0 4
503 321
510 321
510 510
521 510
3 2 11 0 0 4224 0 13 8 0 0 3
927 499
927 478
947 478
3 1 12 0 0 4224 0 14 8 0 0 3
926 438
926 460
947 460
3 2 13 0 0 4224 0 11 9 0 0 3
750 487
750 473
756 473
3 1 14 0 0 4224 0 12 9 0 0 3
750 434
750 455
756 455
3 2 15 0 0 4224 0 15 10 0 0 3
566 501
566 483
584 483
3 1 16 0 0 4224 0 16 10 0 0 3
566 446
566 465
584 465
0 0 17 0 0 4096 0 0 0 24 18 2
503 492
503 538
0 0 17 0 0 4096 0 0 0 23 18 2
693 479
693 538
1 0 17 0 0 4224 0 1 0 0 19 3
414 538
873 538
873 490
1 1 17 0 0 0 0 5 13 0 0 3
864 487
864 490
882 490
2 2 18 0 0 8320 0 5 14 0 0 3
864 451
864 447
881 447
2 2 19 0 0 4224 0 6 12 0 0 2
682 443
705 443
2 2 20 0 0 4224 0 7 16 0 0 2
492 455
521 455
1 1 17 0 0 0 0 6 11 0 0 3
682 479
705 479
705 478
1 1 17 0 0 0 0 7 15 0 0 3
492 491
492 492
521 492
1 0 21 0 0 4096 0 32 0 0 33 2
1084 305
1084 304
1 0 6 0 0 0 0 31 0 0 35 2
713 303
713 302
1 0 5 0 0 0 0 30 0 0 34 2
894 302
894 301
1 0 7 0 0 0 0 29 0 0 36 2
528 303
528 303
0 1 7 0 0 128 0 0 22 36 0 4
506 303
506 188
464 188
464 157
0 2 6 0 0 8320 0 0 22 35 0 4
694 302
694 184
458 184
458 157
0 3 5 0 0 8320 0 0 22 34 0 4
871 301
871 178
452 178
452 157
0 4 21 0 0 8320 0 0 22 33 0 4
1064 304
1064 172
446 172
446 157
6 1 21 0 0 0 0 20 27 0 0 3
1055 303
1055 304
1121 304
6 1 5 0 0 0 0 19 26 0 0 2
857 301
928 301
6 1 6 0 0 0 0 18 25 0 0 2
687 302
744 302
6 1 7 0 0 0 0 17 24 0 0 2
497 303
564 303
1 2 22 0 0 4224 0 23 17 0 0 4
364 308
437 308
437 312
442 312
1 1 22 0 0 0 0 28 23 0 0 3
353 357
353 308
364 308
3 2 23 0 0 8320 0 21 28 0 0 3
314 306
319 306
319 353
1 3 22 0 0 4224 24 4 28 0 0 2
321 361
319 361
4 0 25 0 0 4096 0 17 0 0 44 2
473 351
473 363
4 0 25 0 0 4096 0 18 0 0 44 2
663 350
663 363
4 0 25 0 0 4096 0 19 0 0 44 2
833 349
833 363
1 4 25 0 0 4224 0 3 20 0 0 3
421 363
1031 363
1031 351
1 0 26 0 0 4096 0 17 0 0 46 2
449 303
427 303
0 3 26 0 0 4096 0 0 17 52 0 3
427 209
427 321
449 321
1 0 26 0 0 0 0 18 0 0 48 2
639 302
622 302
0 3 26 0 0 0 0 0 18 52 0 3
622 209
622 320
639 320
1 0 26 0 0 0 0 19 0 0 50 2
809 301
793 301
0 3 26 0 0 0 0 0 19 52 0 3
793 209
793 319
809 319
1 0 26 0 0 0 0 20 0 0 52 2
1007 303
983 303
1 3 26 0 0 4224 0 2 20 0 0 4
312 209
983 209
983 321
1007 321
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
