CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 636 1536 824
193986578 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 275 263 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 375 265 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 266 111 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
14 Logic Display~
6 1050 189 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 679 187 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 860 186 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 494 187 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
12 SPDT Switch~
164 302 259 0 10 11
0 6 6 8 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3747 0 0
0
0
5 SCOPE
12 1087 194 0 1 11
0 2
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 894 191 0 1 11
0 4
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 710 192 0 1 11
0 3
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9325 0 0
0
0
5 SCOPE
12 530 193 0 1 11
0 5
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8903 0 0
0
0
5 SCOPE
12 330 198 0 1 11
0 6
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3834 0 0
0
0
12 Hex Display~
7 421 35 0 18 19
10 5 3 4 2 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3363 0 0
0
0
7 Pulser~
4 256 217 0 10 12
0 11 12 6 13 0 0 5 5 4
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7668 0 0
0
0
6 JK RN~
219 997 222 0 6 22
0 10 4 10 9 14 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 2 0
1 U
4718 0 0
0
0
6 JK RN~
219 799 220 0 6 22
0 10 3 10 9 15 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 2 0
1 U
3874 0 0
0
0
6 JK RN~
219 629 221 0 6 22
0 10 5 10 9 16 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 2 1 0
1 U
6671 0 0
0
0
6 JK RN~
219 439 222 0 6 22
0 10 6 10 9 17 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 512 2 1 1 0
1 U
3789 0 0
0
0
31
1 0 2 0 0 4096 0 4 0 0 9 2
1050 207
1050 206
1 0 3 0 0 4096 0 5 0 0 11 2
679 205
679 204
1 0 4 0 0 4096 0 6 0 0 10 2
860 204
860 203
1 0 5 0 0 0 0 7 0 0 12 2
494 205
494 205
0 1 5 0 0 4224 0 0 14 12 0 4
472 205
472 90
430 90
430 59
0 2 3 0 0 8320 0 0 14 11 0 4
660 204
660 86
424 86
424 59
0 3 4 0 0 8336 0 0 14 10 0 4
837 203
837 80
418 80
418 59
0 4 2 0 0 8320 0 0 14 9 0 4
1030 206
1030 74
412 74
412 59
6 1 2 0 0 0 0 16 9 0 0 3
1021 205
1021 206
1087 206
6 1 4 0 0 0 0 17 10 0 0 2
823 203
894 203
6 1 3 0 0 0 0 18 11 0 0 2
653 204
710 204
6 1 5 0 0 0 0 19 12 0 0 2
463 205
530 205
2 1 4 0 0 0 0 16 10 0 0 3
966 214
894 214
894 203
2 1 5 0 0 0 0 18 12 0 0 3
598 213
530 213
530 205
2 1 3 0 0 0 0 17 11 0 0 3
768 212
710 212
710 204
1 2 6 0 0 4224 0 13 19 0 0 4
330 210
403 210
403 214
408 214
1 1 6 0 0 0 0 8 13 0 0 3
319 259
319 210
330 210
3 2 6 0 0 8320 7 15 8 0 0 3
280 208
285 208
285 255
1 3 8 0 0 4224 0 1 8 0 0 2
287 263
285 263
4 0 9 0 0 4096 0 19 0 0 23 2
439 253
439 265
4 0 9 0 0 4096 0 18 0 0 23 2
629 252
629 265
4 0 9 0 0 4096 0 17 0 0 23 2
799 251
799 265
1 4 9 0 0 4224 0 2 16 0 0 3
387 265
997 265
997 253
1 0 10 0 0 4096 0 19 0 0 25 2
415 205
393 205
0 3 10 0 0 4096 0 0 19 31 0 3
393 111
393 223
415 223
1 0 10 0 0 0 0 18 0 0 27 2
605 204
588 204
0 3 10 0 0 0 0 0 18 31 0 3
588 111
588 222
605 222
1 0 10 0 0 0 0 17 0 0 29 2
775 203
759 203
0 3 10 0 0 0 0 0 17 31 0 3
759 111
759 221
775 221
1 0 10 0 0 0 0 16 0 0 31 2
973 205
949 205
1 3 10 0 0 4224 0 3 16 0 0 4
278 111
949 111
949 223
973 223
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
