CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 830 30 100 9
769 79 1535 823
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
769 79 1535 823
177209362 0
0
6 Title:
5 Name:
0
0
0
41
13 Logic Switch~
5 335 1170 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 333 1111 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 279 1262 0 1 11
0 2
0
0 0 21360 90
2 0V
14 0 28 8
3 V15
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 55 1056 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 58 964 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 161 858 0 1 11
0 15
0
0 0 21360 90
2 0V
14 0 28 8
3 V12
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 51 767 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 55 657 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 61 539 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 61 481 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 62 440 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 63 391 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 63 338 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 66 291 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3363 0 0
0
0
13 Logic Switch~
5 65 247 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7668 0 0
0
0
13 Logic Switch~
5 66 200 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4718 0 0
0
0
13 Logic Switch~
5 65 159 0 1 11
0 38
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3874 0 0
0
0
14 Logic Display~
6 658 1081 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
8 2-In OR~
219 564 1123 0 3 22
0 5 6 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3789 0 0
0
0
9 2-In AND~
219 486 1171 0 3 22
0 2 8 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
4871 0 0
0
0
9 2-In AND~
219 499 1075 0 3 22
0 9 7 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3750 0 0
0
0
9 Inverter~
13 413 1134 0 2 22
0 2 7
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
8778 0 0
0
0
14 Logic Display~
6 374 959 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
538 0 0
0
0
8 2-In OR~
219 282 995 0 3 22
0 12 11 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6843 0 0
0
0
9 2-In AND~
219 210 1041 0 3 22
0 2 14 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3136 0 0
0
0
9 2-In AND~
219 212 960 0 3 22
0 13 3 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
5950 0 0
0
0
9 Inverter~
13 116 1009 0 2 22
0 2 3
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U2F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
5670 0 0
0
0
14 Logic Display~
6 366 667 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6828 0 0
0
0
8 2-In OR~
219 289 702 0 3 22
0 17 18 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6735 0 0
0
0
9 2-In AND~
219 213 743 0 3 22
0 15 19 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8365 0 0
0
0
9 2-In AND~
219 215 654 0 3 22
0 20 21 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4132 0 0
0
0
9 Inverter~
13 130 706 0 2 22
0 15 21
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U2E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
4551 0 0
0
0
14 Logic Display~
6 466 297 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3635 0 0
0
0
14 Logic Display~
6 463 253 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3973 0 0
0
0
14 Logic Display~
6 456 206 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3851 0 0
0
0
14 Logic Display~
6 440 150 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8383 0 0
0
0
9 Inverter~
13 385 265 0 2 22
0 26 22
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9334 0 0
0
0
9 Inverter~
13 351 246 0 2 22
0 27 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
7471 0 0
0
0
9 Inverter~
13 371 228 0 2 22
0 28 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3334 0 0
0
0
9 Inverter~
13 355 207 0 2 22
0 29 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3559 0 0
0
0
5 74147
219 267 241 0 13 27
0 38 37 36 35 34 33 32 31 30
26 27 28 29
0
0 0 13040 0
5 74147
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
121 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
27

0 10 5 4 3 2 1 13 12 11
9 7 6 14 10 5 4 3 2 1
13 12 11 9 7 6 14 0
65 0 0 0 1 0 0 0
1 U
984 0 0
0
0
41
1 0 2 0 0 8192 0 3 0 0 8 4
280 1249
280 1159
438 1159
438 1162
0 1 2 0 0 4224 0 0 3 4 0 4
152 1032
152 1242
280 1242
280 1249
2 2 3 0 0 4224 0 26 27 0 0 3
188 969
119 969
119 991
1 1 2 0 0 0 0 27 25 0 0 3
119 1027
119 1032
186 1032
3 1 4 0 0 4224 0 19 18 0 0 3
597 1123
658 1123
658 1099
1 3 5 0 0 8320 0 19 21 0 0 4
551 1114
528 1114
528 1075
520 1075
3 2 6 0 0 8320 0 20 19 0 0 4
507 1171
543 1171
543 1132
551 1132
1 1 2 0 0 0 0 20 22 0 0 3
462 1162
416 1162
416 1152
2 2 7 0 0 8320 0 22 21 0 0 3
416 1116
416 1084
475 1084
2 1 8 0 0 4224 0 20 1 0 0 4
462 1180
356 1180
356 1170
347 1170
1 1 9 0 0 4224 0 2 21 0 0 4
345 1111
467 1111
467 1066
475 1066
3 1 10 0 0 4224 0 24 23 0 0 3
315 995
374 995
374 977
2 3 11 0 0 8320 0 24 25 0 0 4
269 1004
239 1004
239 1041
231 1041
3 1 12 0 0 4224 0 26 24 0 0 4
233 960
261 960
261 986
269 986
1 1 13 0 0 4224 0 5 26 0 0 4
70 964
180 964
180 951
188 951
1 2 14 0 0 4224 0 4 25 0 0 4
67 1056
178 1056
178 1050
186 1050
0 1 15 0 0 4224 0 0 6 24 0 4
163 734
163 838
162 838
162 845
3 1 16 0 0 4224 0 29 28 0 0 3
322 702
366 702
366 685
1 3 17 0 0 8320 0 29 31 0 0 4
276 693
244 693
244 654
236 654
3 2 18 0 0 4224 0 30 29 0 0 4
234 743
268 743
268 711
276 711
1 2 19 0 0 4224 0 7 30 0 0 4
63 767
181 767
181 752
189 752
1 1 20 0 0 4224 0 8 31 0 0 4
67 657
183 657
183 645
191 645
2 2 21 0 0 8320 0 32 31 0 0 3
133 688
133 663
191 663
1 1 15 0 0 0 0 30 32 0 0 3
189 734
133 734
133 724
2 1 22 0 0 8336 0 37 33 0 0 5
406 265
425 265
425 321
466 321
466 315
1 2 23 0 0 8320 0 34 38 0 0 4
463 271
463 269
372 269
372 246
1 2 24 0 0 8320 0 35 39 0 0 3
456 224
456 228
392 228
2 1 25 0 0 4224 0 40 36 0 0 3
376 207
440 207
440 168
1 10 26 0 0 4224 0 37 41 0 0 4
370 265
313 265
313 250
305 250
11 1 27 0 0 4224 0 41 38 0 0 4
305 241
328 241
328 246
336 246
1 12 28 0 0 4224 0 39 41 0 0 4
356 228
313 228
313 232
305 232
13 1 29 0 0 4224 0 41 40 0 0 4
305 223
332 223
332 207
340 207
1 9 30 0 0 8320 0 9 41 0 0 4
73 539
221 539
221 277
229 277
8 1 31 0 0 8320 0 41 10 0 0 4
229 268
84 268
84 481
73 481
1 7 32 0 0 8320 0 11 41 0 0 4
74 440
221 440
221 259
229 259
6 1 33 0 0 4224 0 41 12 0 0 4
229 250
84 250
84 391
75 391
1 5 34 0 0 4224 0 13 41 0 0 4
75 338
221 338
221 241
229 241
4 1 35 0 0 4224 0 41 14 0 0 4
229 232
87 232
87 291
78 291
1 3 36 0 0 4224 0 15 41 0 0 4
77 247
221 247
221 223
229 223
2 1 37 0 0 4224 0 41 16 0 0 4
229 214
87 214
87 200
78 200
1 1 38 0 0 4224 0 17 41 0 0 4
77 159
221 159
221 205
229 205
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
