CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
769 79 2305 832
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
769 79 2305 832
177209362 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 315 433 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 70 436 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 349 369 0 1 11
0 8
0
0 0 21360 90
2 0V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 315 369 0 1 11
0 9
0
0 0 21360 90
2 0V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 150 368 0 1 11
0 6
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 118 366 0 1 11
0 7
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
14 Logic Display~
6 378 255 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 361 254 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 343 256 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 325 253 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 181 250 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 163 253 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 144 251 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 126 252 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
6 74LS90
107 352 308 0 10 21
0 9 9 8 8 3 4 3 12 11
10
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U2
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
6 74LS90
107 153 304 0 10 21
0 7 7 6 6 5 2 15 14 13
2
0
0 0 13040 90
6 74LS90
-21 -51 21 -43
2 U1
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
20
1 6 2 0 0 4224 0 11 16 0 0 3
181 268
181 336
180 336
5 1 3 0 0 12416 0 15 10 0 0 6
370 340
370 344
306 344
306 237
325 237
325 271
6 1 4 0 0 4224 0 15 1 0 0 3
379 340
379 433
327 433
5 1 5 0 0 4224 0 16 2 0 0 3
171 336
171 436
82 436
4 0 6 0 0 4096 0 16 0 0 11 4
153 330
153 343
151 343
151 348
1 2 7 0 0 8320 0 6 16 0 0 4
119 353
119 344
135 344
135 330
1 4 8 0 0 12288 0 3 15 0 0 4
350 356
350 348
352 348
352 334
3 1 8 0 0 4224 0 15 3 0 0 4
343 334
343 349
350 349
350 356
2 1 9 0 0 8320 0 15 4 0 0 4
334 334
334 349
316 349
316 356
1 1 9 0 0 0 0 15 4 0 0 4
325 334
325 349
316 349
316 356
3 1 6 0 0 4224 0 16 5 0 0 4
144 330
144 348
151 348
151 355
1 1 7 0 0 0 0 6 16 0 0 4
119 353
119 344
126 344
126 330
1 10 10 0 0 4224 0 7 15 0 0 3
378 273
378 270
379 270
1 9 11 0 0 4224 0 8 15 0 0 2
361 272
361 270
1 8 12 0 0 4224 0 9 15 0 0 2
343 274
343 270
1 7 3 0 0 0 0 10 15 0 0 2
325 271
325 270
1 10 2 0 0 0 0 11 16 0 0 3
181 268
181 266
180 266
1 9 13 0 0 4224 0 12 16 0 0 3
163 271
163 266
162 266
1 8 14 0 0 4224 0 13 16 0 0 2
144 269
144 266
1 7 15 0 0 4224 0 14 16 0 0 2
126 270
126 266
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
