CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 890 30 100 9
769 79 1535 823
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
769 79 1535 823
177209362 0
0
6 Title:
5 Name:
0
0
0
39
13 Logic Switch~
5 194 936 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 195 895 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 194 847 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 194 802 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 131 784 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 165 538 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 31 483 0 1 11
0 16
0
0 0 21360 0
2 0V
-8 -17 6 -9
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 29 449 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 30 410 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 30 365 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 23 207 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 25 143 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 43 43 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3834 0 0
0
0
9 CA 7-Seg~
184 235 621 0 18 19
10 13 12 11 10 9 8 7 39 14
0 0 0 0 0 0 0 2 1
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3363 0 0
0
0
6 74LS47
187 230 729 0 14 29
0 2 3 4 5 6 40 7 8 9
10 11 12 13 41
0
0 0 13040 602
6 74LS47
-21 -60 21 -52
2 U4
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7668 0 0
0
0
14 Logic Display~
6 518 331 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 495 333 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 462 332 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 427 333 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 393 329 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 363 330 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 336 331 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 309 333 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 285 333 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
14 Logic Display~
6 262 334 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3136 0 0
0
0
6 74LS42
101 165 406 0 14 29
0 28 27 15 16 17 18 19 20 21
22 23 24 25 26
0
0 0 13040 0
6 74LS42
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 11 10 9 7 6
5 4 3 2 1 12 13 14 15 11
10 9 7 6 5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
5950 0 0
0
0
14 Logic Display~
6 448 263 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5670 0 0
0
0
14 Logic Display~
6 440 221 0 1 2
10 36
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6828 0 0
0
0
14 Logic Display~
6 439 175 0 1 2
10 35
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6735 0 0
0
0
14 Logic Display~
6 435 118 0 1 2
10 34
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8365 0 0
0
0
10 2-In NAND~
219 382 285 0 3 22
0 30 29 37
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
4132 0 0
0
0
10 2-In NAND~
219 383 246 0 3 22
0 29 33 36
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4551 0 0
0
0
10 2-In NAND~
219 382 198 0 3 22
0 30 31 35
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3635 0 0
0
0
10 2-In NAND~
219 381 150 0 3 22
0 33 31 34
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3973 0 0
0
0
9 Inverter~
13 125 207 0 2 22
0 29 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3851 0 0
0
0
9 Inverter~
13 170 141 0 2 22
0 30 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8383 0 0
0
0
14 Logic Display~
6 207 60 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9334 0 0
0
0
14 Logic Display~
6 207 15 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7471 0 0
0
0
9 Inverter~
13 133 43 0 2 22
0 32 38
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3334 0 0
0
0
55
1 1 2 0 0 4224 0 15 1 0 0 3
271 766
271 936
206 936
1 2 3 0 0 8320 0 2 15 0 0 3
207 895
262 895
262 766
3 1 4 0 0 4224 0 15 3 0 0 3
253 766
253 847
206 847
4 1 5 0 0 8320 0 15 4 0 0 3
244 766
244 802
206 802
1 5 6 0 0 4224 0 5 15 0 0 3
143 784
199 784
199 766
7 7 7 0 0 4224 0 15 14 0 0 4
271 696
271 665
250 665
250 657
6 8 8 0 0 4224 0 14 15 0 0 4
244 657
244 688
262 688
262 696
9 5 9 0 0 4224 0 15 14 0 0 4
253 696
253 665
238 665
238 657
4 10 10 0 0 4224 0 14 15 0 0 4
232 657
232 688
244 688
244 696
11 3 11 0 0 4224 0 15 14 0 0 4
235 696
235 665
226 665
226 657
2 12 12 0 0 4224 0 14 15 0 0 4
220 657
220 688
226 688
226 696
13 1 13 0 0 4224 0 15 14 0 0 4
217 696
217 665
214 665
214 657
1 9 14 0 0 4224 0 6 14 0 0 3
177 538
235 538
235 585
1 3 15 0 0 4224 0 8 26 0 0 4
41 449
125 449
125 442
133 442
1 4 16 0 0 4224 0 7 26 0 0 4
43 483
125 483
125 451
133 451
1 9 17 0 0 4096 0 16 0 0 36 3
518 349
518 359
519 359
1 8 18 0 0 4096 0 17 0 0 36 2
495 351
495 359
1 7 19 0 0 4096 0 18 0 0 36 3
462 350
462 359
464 359
1 6 20 0 0 4096 0 19 0 0 36 2
427 351
427 359
1 5 21 0 0 4224 0 20 0 0 36 2
393 347
393 359
1 4 22 0 0 4096 0 21 0 0 36 2
363 348
363 359
1 3 23 0 0 4096 0 22 0 0 36 2
336 349
336 359
1 2 24 0 0 4096 0 23 0 0 36 3
309 351
309 359
311 359
1 1 25 0 0 4096 0 24 0 0 36 3
285 351
285 359
283 359
1 0 26 0 0 4096 0 25 0 0 36 3
262 352
262 359
259 359
5 9 17 0 0 4224 0 26 0 0 36 2
203 370
217 370
6 8 18 0 0 4224 0 26 0 0 36 2
203 379
217 379
7 7 19 0 0 4224 0 26 0 0 36 2
203 388
217 388
8 6 20 0 0 4224 0 26 0 0 36 2
203 397
217 397
9 5 21 0 0 0 0 26 0 0 36 4
203 406
212 406
212 407
217 407
10 4 22 0 0 4224 0 26 0 0 36 2
203 415
217 415
11 3 23 0 0 4224 0 26 0 0 36 2
203 424
217 424
12 2 24 0 0 4224 0 26 0 0 36 2
203 433
217 433
13 1 25 0 0 4224 0 26 0 0 36 2
203 442
217 442
14 0 26 0 0 4224 0 26 0 0 36 2
203 451
217 451
10 0 1 0 0 8352 0 0 0 0 0 3
217 462
217 359
535 359
1 2 27 0 0 4224 0 9 26 0 0 4
42 410
125 410
125 433
133 433
1 1 28 0 0 4224 0 10 26 0 0 4
42 365
125 365
125 424
133 424
0 2 29 0 0 8320 0 0 31 45 0 3
69 207
69 294
358 294
0 1 30 0 0 8320 0 0 31 46 0 3
86 141
86 276
358 276
0 1 29 0 0 0 0 0 32 45 0 3
96 207
96 237
359 237
0 1 30 0 0 0 0 0 33 46 0 3
144 141
144 189
358 189
0 2 31 0 0 8192 0 0 34 44 0 3
307 207
307 159
357 159
2 2 31 0 0 4240 0 35 33 0 0 2
146 207
358 207
1 1 29 0 0 0 0 11 35 0 0 2
35 207
110 207
1 1 30 0 0 0 0 12 36 0 0 3
37 143
37 141
155 141
1 0 32 0 0 8320 0 37 0 0 55 4
207 78
207 86
97 86
97 43
2 0 33 0 0 8192 0 32 0 0 49 3
359 255
298 255
298 141
2 1 33 0 0 4224 0 36 34 0 0 2
191 141
357 141
1 3 34 0 0 8320 0 30 34 0 0 3
435 136
435 150
408 150
3 1 35 0 0 4224 0 33 29 0 0 3
409 198
439 198
439 193
1 3 36 0 0 8320 0 28 32 0 0 3
440 239
440 246
410 246
3 1 37 0 0 4224 0 31 27 0 0 3
409 285
448 285
448 281
1 2 38 0 0 8320 0 38 39 0 0 3
207 33
207 43
154 43
1 1 32 0 0 0 0 13 39 0 0 2
55 43
118 43
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
