CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
42991634 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 217 199 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 97 271 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
14 Logic Display~
6 807 120 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
5 SCOPE
12 834 125 0 1 11
0 2
0
0 0 57584 0
3 TP6
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6153 0 0
0
0
9 Inverter~
13 188 141 0 2 22
0 3 4
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
5394 0 0
0
0
5 SCOPE
12 684 125 0 1 11
0 5
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 517 125 0 1 11
0 6
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 341 126 0 1 11
0 7
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 207 228 0 1 11
0 8
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3549 0 0
0
0
14 Logic Display~
6 651 117 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 484 119 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 315 118 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
6 JK RN~
219 269 153 0 6 22
0 3 8 4 14 13 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 1 0
1 U
3834 0 0
0
0
6 JK RN~
219 439 153 0 6 22
0 7 8 13 14 12 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 1 0
1 U
3363 0 0
0
0
6 JK RN~
219 611 153 0 6 22
0 6 8 12 14 11 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 2 0
1 U
7668 0 0
0
0
6 JK RN~
219 768 153 0 6 22
0 5 8 11 14 3 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 2 0
1 U
4718 0 0
0
0
12 SPDT Switch~
164 167 239 0 10 11
0 8 8 9 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3874 0 0
0
0
7 Pulser~
4 91 207 0 10 12
0 15 16 8 17 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6671 0 0
0
0
28
1 0 2 0 0 4096 0 3 0 0 3 2
807 138
807 137
5 0 3 0 0 12432 0 16 0 0 5 5
798 154
894 154
894 74
215 74
215 119
6 1 2 0 0 8320 0 16 4 0 0 3
792 136
792 137
834 137
2 3 4 0 0 8320 0 5 13 0 0 5
191 159
191 163
230 163
230 154
245 154
1 1 3 0 0 0 0 5 13 0 0 5
191 123
191 119
230 119
230 136
245 136
1 0 5 0 0 4096 0 6 0 0 20 2
684 137
684 136
1 0 6 0 0 4096 0 7 0 0 22 2
517 137
517 136
1 0 7 0 0 4096 0 8 0 0 24 2
341 138
341 136
1 0 8 0 0 4096 0 9 0 0 16 2
207 240
207 239
1 0 5 0 0 0 0 10 0 0 20 2
651 135
651 136
1 0 6 0 0 0 0 11 0 0 22 2
484 137
484 136
1 0 7 0 0 0 0 12 0 0 24 2
315 136
315 136
0 2 8 0 0 4096 0 0 16 14 0 4
572 237
729 237
729 145
737 145
0 2 8 0 0 4224 0 0 15 15 0 4
390 237
572 237
572 145
580 145
2 0 8 0 0 0 0 14 0 0 16 5
408 145
390 145
390 238
233 238
233 239
1 2 8 0 0 0 0 17 13 0 0 4
184 239
235 239
235 145
238 145
3 1 9 0 0 4224 0 17 2 0 0 4
150 243
118 243
118 271
109 271
3 2 8 0 0 8320 10 18 17 0 0 4
115 198
142 198
142 235
150 235
5 3 11 0 0 4224 0 15 16 0 0 2
641 154
744 154
6 1 5 0 0 4224 0 15 16 0 0 2
635 136
744 136
5 3 12 0 0 4224 0 14 15 0 0 2
469 154
587 154
6 1 6 0 0 4224 0 14 15 0 0 2
463 136
587 136
5 3 13 0 0 4224 0 13 14 0 0 2
299 154
415 154
6 1 7 0 0 4224 0 13 14 0 0 2
293 136
415 136
4 0 14 0 0 8192 0 16 0 0 26 3
768 184
768 197
611 197
4 0 14 0 0 8320 0 15 0 0 27 4
611 184
611 197
438 197
438 198
0 4 14 0 0 0 0 0 14 28 0 4
268 199
268 198
439 198
439 184
1 4 14 0 0 0 0 1 13 0 0 3
229 199
269 199
269 184
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
